import video_modes_pkg::*;
import clock_modes_pkg::*;

module Top (
    // Fun stuff
    input logic btn,
    output logic led,
    output logic [7:0] seg,

    // Borin stuff
    input logic clk_ext, // 100MHz for now
    input logic reset,

    // SPI (Slave)
    input logic spi_sclk,
    input logic spi_ssn,
    input logic spi_mosi,
    output logic spi_miso,

    // VGA control
    output logic vga_hsync,
    output logic vga_vsync,
    output logic[3:0] vga_red,
    output logic[3:0] vga_green,
    output logic[3:0] vga_blue
);
    localparam video_mode_t VIDEO_MODE = VMODE_640x480p60;

    assign led = btn;

    ////////////////////////////////////////////////
    ////////////// CLOCK GENERATION ////////////////
    ////////////////////////////////////////////////

    logic clk_display;
    logic rstn_display;

    logic clk_system;
    logic rstn_system;

    ClockManager #(
        .CLK_DISPLAY(VIDEO_MODE.clock_config),
        .CLK_SYSTEM(CLK_100_50_MHZ)
    ) clock_manager_inst (
        .clk_ext(clk_ext),
        .reset(reset),

        .clk_system(clk_system),
        .rstn_system(rstn_system),

        .clk_display(clk_display),
        .rstn_display(rstn_display)
    );


    ///////////////////////////////////////
    ////////////// DISPLAY ////////////////
    ///////////////////////////////////////

    Display #(
        .VIDEO_MODE(VIDEO_MODE)
    ) display_inst (
        .clk_pixel(clk_display),
        .rstn_pixel(rstn_display),

        .vga_hsync(vga_hsync),
        .vga_vsync(vga_vsync),
        .vga_red(vga_red),
        .vga_green(vga_green),
        .vga_blue(vga_blue)
    );

    logic [7:0] spi_data_rx;
    logic spi_data_ready;

    Spi spi_inst (
        .sclk(spi_sclk),
        .ssn(spi_ssn),
        .miso(spi_miso),
        .mosi(spi_mosi),
        .data_rx(spi_data_rx),
        .data_ready(spi_data_ready)
    );

    always_ff @(posedge clk_system or negedge rstn_system) begin
        if (!rstn_system) begin
            seg <= 8'b0;
        end else begin
            if (spi_data_ready) begin
                seg <= ~spi_data_rx;
            end
        end
    end

endmodule


