package reciprocal_divider_params;
    // MUST MATCH THE DIVIDER XCI FILE!
    parameter int DIVIDEND_AND_QUOTIENT_WIDTH = 56; // Ops, this one is always 6 above for some reason.
    parameter int DIVISOR_WIDTH = 32;
    parameter int DIVIDER_LATENCY = 10;
endpackage
