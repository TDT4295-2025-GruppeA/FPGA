module PipelineTail();


    

endmodule