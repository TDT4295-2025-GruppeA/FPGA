// Example module used to demonstrate the test system
// Simply adds two integers
module Example(
    input int a,
    input int b,
    output int sum
);
    assign sum = a + b;
endmodule
