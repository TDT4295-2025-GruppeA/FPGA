import fixed_pkg::*;

package types_pkg;
    typedef struct packed {
        logic [3:0] red;
        logic [3:0] green;
        logic [3:0] blue;
    } color_t;

    typedef struct packed {
        fixed x;
        fixed y;
        fixed z;
    } position_t;

    typedef struct packed {
        position_t position;
        color_t color;
    } vertex_t;

    typedef struct packed {
        vertex_t v0;
        vertex_t v1;
        vertex_t v2;
    } triangle_t;

    typedef struct packed {
        fixed m00;
        fixed m01;
        fixed m02;
        fixed m10;
        fixed m11;
        fixed m12;
        fixed m20;
        fixed m21;
        fixed m22;
    } rotmat_t;

    typedef struct packed {
        position_t position;
        rotmat_t rotmat;
    } transform_t;

    typedef struct packed {
        logic [7:0] model_id;
        transform_t transform;
    } modelinstance_t;

    typedef struct packed {
        triangle_t triangle;
        transform_t transform;
    } triangle_tf_t;

endpackage