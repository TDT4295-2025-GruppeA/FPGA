

module Top (
    input btn[4],
    output led[4]
);
    assign led = btn;

endmodule;


